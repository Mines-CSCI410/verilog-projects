module student_half_adder(input a, b, output sum, carry);
    // Details in the textbook.
endmodule
