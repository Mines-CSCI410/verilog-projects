module student_add16(input [15:0] a, b, output [15:0] out);
    // Implement a 16 bit adder (without using assign out = a + b)
endmodule
