module student_alu(
    // Implement an ALU here, details are in the textbook.
endmodule
