module student_full_adder(input a, b, c, output sum, carry);
    // Details in the textbook.
endmodule
