module student_bit (input in, load, output out);
endmodule
