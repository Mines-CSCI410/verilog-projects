module mux8way16_test;
  reg [15:0] a, b, c, d, e, f, g, h;
  reg [2:0] sel;
  wire [15:0] out;

  student_mux8way16 dut (.a(a), .b(b), .c(c), .d(d), .e(e), .f(f), .g(g), .h(h), .sel(sel), .out(out));

  initial begin
    $display("|a|b|c|d|e|f|g|h|sel|out|");

    a = 'b0000000000000000;
    b = 'b0000000000000000;
    c = 'b0000000000000000;
    d = 'b0000000000000000;
    e = 'b0000000000000000;
    f = 'b0000000000000000;
    g = 'b0000000000000000;
    h = 'b0000000000000000;
    sel = 'b000;
    #1 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0000000000000000;
    b = 'b0000000000000000;
    c = 'b0000000000000000;
    d = 'b0000000000000000;
    e = 'b0000000000000000;
    f = 'b0000000000000000;
    g = 'b0000000000000000;
    h = 'b0000000000000000;
    sel = 'b001;
    #2 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0000000000000000;
    b = 'b0000000000000000;
    c = 'b0000000000000000;
    d = 'b0000000000000000;
    e = 'b0000000000000000;
    f = 'b0000000000000000;
    g = 'b0000000000000000;
    h = 'b0000000000000000;
    sel = 'b010;
    #3 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0000000000000000;
    b = 'b0000000000000000;
    c = 'b0000000000000000;
    d = 'b0000000000000000;
    e = 'b0000000000000000;
    f = 'b0000000000000000;
    g = 'b0000000000000000;
    h = 'b0000000000000000;
    sel = 'b011;
    #4 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0000000000000000;
    b = 'b0000000000000000;
    c = 'b0000000000000000;
    d = 'b0000000000000000;
    e = 'b0000000000000000;
    f = 'b0000000000000000;
    g = 'b0000000000000000;
    h = 'b0000000000000000;
    sel = 'b100;
    #5 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0000000000000000;
    b = 'b0000000000000000;
    c = 'b0000000000000000;
    d = 'b0000000000000000;
    e = 'b0000000000000000;
    f = 'b0000000000000000;
    g = 'b0000000000000000;
    h = 'b0000000000000000;
    sel = 'b101;
    #6 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0000000000000000;
    b = 'b0000000000000000;
    c = 'b0000000000000000;
    d = 'b0000000000000000;
    e = 'b0000000000000000;
    f = 'b0000000000000000;
    g = 'b0000000000000000;
    h = 'b0000000000000000;
    sel = 'b110;
    #7 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0000000000000000;
    b = 'b0000000000000000;
    c = 'b0000000000000000;
    d = 'b0000000000000000;
    e = 'b0000000000000000;
    f = 'b0000000000000000;
    g = 'b0000000000000000;
    h = 'b0000000000000000;
    sel = 'b111;
    #8 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0001001000110100;
    b = 'b0010001101000101;
    c = 'b0011010001010110;
    d = 'b0100010101100111;
    e = 'b0101011001111000;
    f = 'b0110011110001001;
    g = 'b0111100010011010;
    h = 'b1000100110101011;
    sel = 'b000;
    #9 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0001001000110100;
    b = 'b0010001101000101;
    c = 'b0011010001010110;
    d = 'b0100010101100111;
    e = 'b0101011001111000;
    f = 'b0110011110001001;
    g = 'b0111100010011010;
    h = 'b1000100110101011;
    sel = 'b001;
    #10 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0001001000110100;
    b = 'b0010001101000101;
    c = 'b0011010001010110;
    d = 'b0100010101100111;
    e = 'b0101011001111000;
    f = 'b0110011110001001;
    g = 'b0111100010011010;
    h = 'b1000100110101011;
    sel = 'b010;
    #11 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0001001000110100;
    b = 'b0010001101000101;
    c = 'b0011010001010110;
    d = 'b0100010101100111;
    e = 'b0101011001111000;
    f = 'b0110011110001001;
    g = 'b0111100010011010;
    h = 'b1000100110101011;
    sel = 'b011;
    #12 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0001001000110100;
    b = 'b0010001101000101;
    c = 'b0011010001010110;
    d = 'b0100010101100111;
    e = 'b0101011001111000;
    f = 'b0110011110001001;
    g = 'b0111100010011010;
    h = 'b1000100110101011;
    sel = 'b100;
    #13 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0001001000110100;
    b = 'b0010001101000101;
    c = 'b0011010001010110;
    d = 'b0100010101100111;
    e = 'b0101011001111000;
    f = 'b0110011110001001;
    g = 'b0111100010011010;
    h = 'b1000100110101011;
    sel = 'b101;
    #14 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0001001000110100;
    b = 'b0010001101000101;
    c = 'b0011010001010110;
    d = 'b0100010101100111;
    e = 'b0101011001111000;
    f = 'b0110011110001001;
    g = 'b0111100010011010;
    h = 'b1000100110101011;
    sel = 'b110;
    #15 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

    a = 'b0001001000110100;
    b = 'b0010001101000101;
    c = 'b0011010001010110;
    d = 'b0100010101100111;
    e = 'b0101011001111000;
    f = 'b0110011110001001;
    g = 'b0111100010011010;
    h = 'b1000100110101011;
    sel = 'b111;
    #16 $display("|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|", a, b, c, d, e, f, g, h, sel, out);

  $finish;
  end
endmodule
