module student_pc (input [15:0] in, input reset, load, inc, output [15:0] out);
endmodule
